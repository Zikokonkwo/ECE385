module game_text(
    input clk,
    input [3:0] dig0, dig1,
    input [9:0] drawX, drawY,
    output text_on,
  output reg [11:0] text_rgb
);

//Display Fail Region

//Display Level Region


  
endmodule
