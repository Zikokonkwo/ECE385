mdoule collision_detection();
end module
