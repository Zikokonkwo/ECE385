module game_char(
    input clk,  
    input reset,
    output reg [11:0] graph_rgb
);
endmodule
